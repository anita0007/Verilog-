module mux8to1(x,y,z,I,S,Y);
input [2:0]S;
input x,y,z;
output Y;
output reg [7:0]I;
wire A,B;

always @(x,y,z)begin
	if(x==0 & y==0 & z==0)begin
		I[0] = 1;
	end
	else if(x==0 & y ==1 & z==0) begin
		I[2] = 1;
	end
	else if(x==0 & y ==1 & z==1) begin
		I[3] = 1;
	end
	else if(x==1 & y ==0 & z==1) begin
		I[5] = 1;
	end
	else if(x==1 & y ==1 & z==1) begin
		I[7] = 1;
	end
end

mux4to1 m40(I[0],0,I[2],I[3],S[1:0],A);
mux4to1 m41(0,I[5],0,I[7],S[1:0],B);
mux2to1 m20(A,B,S[2],Y);

endmodule

module decoder3(X,Y);
input [2:0] X;
output [7:0] Y;

decoder d0(x[0],x[1],x[2],